# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_io__fill10
  CLASS PAD SPACER ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_fd_io__fill10 0 0 ;
  SIZE 10 BY 350 ;
  SYMMETRY X Y R90 ;
  SITE GF_IO_Site ;
  PIN DVDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal3 ;
        RECT 9 134 10 149 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 9 150 10 165 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 9 166 10 181 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 9 182 10 197 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 9 214 10 229 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 9 118 10 125 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 9 206 10 213 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 9 262 10 269 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 9 270 10 277 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 9 278 10 285 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 9 294 10 301 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 9 334 10 341 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0 334 1 341 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0 294 1 301 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0 278 1 285 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0 270 1 277 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0 262 1 269 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0 214 1 229 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0 206 1 213 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0 182 1 197 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0 166 1 181 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0 150 1 165 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0 134 1 149 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0 118 1 125 ;
    END
  END DVDD
  PIN DVSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal3 ;
        RECT 9 70 10 85 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 9 86 10 101 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 9 102 10 117 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 9 230 10 245 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 9 126 10 133 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 9 198 10 205 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 9 286 10 293 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 9 302 10 309 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 9 326 10 333 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 9 342 10 348.39 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0 342 1 348.39 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0 326 1 333 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0 302 1 309 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0 286 1 293 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0 230 1 245 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0 198 1 205 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0 126 1 133 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0 102 1 117 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0 86 1 101 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0 70 1 85 ;
    END
  END DVSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal3 ;
        RECT 9 254 10 261 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 9 310 10 317 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0 310 1 317 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0 254 1 261 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal3 ;
        RECT 9 246 10 253 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 9 318 10 325 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0 318 1 325 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0 246 1 253 ;
    END
  END VSS
  OBS
    LAYER Metal1 ;
      RECT 0 0 10 350 ;
    LAYER Metal2 ;
      RECT 0 0 10 350 ;
    LAYER Metal3 ;
      POLYGON 10 69.72 8.72 69.72 8.72 85.28 10 85.28 10 85.72 8.72 85.72 8.72 101.28 10 101.28 10 101.72 8.72 101.72 8.72 117.28 10 117.28 10 117.72 8.72 117.72 8.72 125.28 10 125.28 10 125.72 8.72 125.72 8.72 133.28 10 133.28 10 133.72 8.72 133.72 8.72 149.28 10 149.28 10 149.72 8.72 149.72 8.72 165.28 10 165.28 10 165.72 8.72 165.72 8.72 181.28 10 181.28 10 181.72 8.72 181.72 8.72 197.28 10 197.28 10 197.72 8.72 197.72 8.72 205.28 10 205.28 10 205.72 8.72 205.72 8.72 213.28 10 213.28 10 213.72 8.72 213.72 8.72 229.28 10 229.28 10 229.72 8.72 229.72 8.72 245.28 10 245.28 10 245.72 8.72 245.72 8.72 253.28 10 253.28 10 253.72 8.72 253.72 8.72 261.28 10 261.28 10 261.72 8.72 261.72 8.72 269.28 10 269.28 10 269.72 8.72 269.72 8.72 277.28 10 277.28 10 277.72 8.72 277.72 8.72 285.28 10 285.28 10 285.72 8.72 285.72 8.72 293.28 10 293.28 10 293.72 8.72 293.72 8.72 301.28 10 301.28 10 301.72 8.72 301.72 8.72 309.28 10 309.28 10 309.72 8.72 309.72 8.72 317.28 10 317.28 10 317.72 8.72 317.72 8.72 325.28 10 325.28 10 325.72 8.72 325.72 8.72 333.28 10 333.28 10 333.72 8.72 333.72 8.72 341.28 10 341.28 10 341.72 8.72 341.72 8.72 348.67 10 348.67 10 350 0 350 0 348.67 1.28 348.67 1.28 341.72 0 341.72 0 341.28 1.28 341.28 1.28 333.72 0 333.72 0 333.28 1.28 333.28 1.28 325.72 0 325.72 0 325.28 1.28 325.28 1.28 317.72 0 317.72 0 317.28 1.28 317.28 1.28 309.72 0 309.72 0 309.28 1.28 309.28 1.28 301.72 0 301.72 0 301.28 1.28 301.28 1.28 293.72 0 293.72 0 293.28 1.28 293.28 1.28 285.72 0 285.72 0 285.28 1.28 285.28 1.28 277.72 0 277.72 0 277.28 1.28 277.28 1.28 269.72 0 269.72 0 269.28 1.28 269.28 1.28 261.72 0 261.72 0 261.28 1.28 261.28 1.28 253.72 0 253.72 0 253.28 1.28 253.28 1.28 245.72 0 245.72 0 245.28 1.28 245.28 1.28 229.72 0 229.72 0 229.28 1.28 229.28 1.28 213.72 0 213.72 0 213.28 1.28 213.28 1.28 205.72 0 205.72 0 205.28 1.28 205.28 1.28 197.72 0 197.72 0 197.28 1.28 197.28 1.28 181.72 0 181.72 0 181.28 1.28 181.28 1.28 165.72 0 165.72 0 165.28 1.28 165.28 1.28 149.72 0 149.72 0 149.28 1.28 149.28 1.28 133.72 0 133.72 0 133.28 1.28 133.28 1.28 125.72 0 125.72 0 125.28 1.28 125.28 1.28 117.72 0 117.72 0 117.28 1.28 117.28 1.28 101.72 0 101.72 0 101.28 1.28 101.28 1.28 85.72 0 85.72 0 85.28 1.28 85.28 1.28 69.72 0 69.72 0 0 10 0 ;
    LAYER Via1 ;
      RECT 0 0 10 350 ;
    LAYER Via2 ;
      RECT 0 0 10 350 ;
  END

END gf180mcu_fd_io__fill10
