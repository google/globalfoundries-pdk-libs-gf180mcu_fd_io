* Copyright 2022 GlobalFoundries PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.SUBCKT gf180mcu_fd_io__dvss DVDD DVSS VDD
M0 n6 n7 DVDD DVDD pmos_6p0 m=1.0 w=15e-6 l=700e-9 nf=1.0 as=6.6e-12 ad=6.6e-12
+ ps=30.88e-6 pd=30.88e-6 nrd=29.333e-3 nrs=29.333e-3 sa=440e-9 sb=440e-9
+ sd=0.0 dtemp=0.0 par=1
M1 n7 n8 DVDD DVDD pmos_6p0 m=1.0 w=20e-6 l=700e-9 nf=1.0 as=8.8e-12 ad=8.8e-12
+ ps=40.88e-6 pd=40.88e-6 nrd=22e-3 nrs=22e-3 sa=440e-9 sb=440e-9 sd=0.0
+ dtemp=0.0 par=1
M2 n4 n6 DVDD DVDD pmos_6p0 m=1.0 w=120e-6 l=700e-9 nf=2.0 as=52.8e-12 ad=31.2e-12
+ ps=241.76e-6 pd=121.04e-6 nrd=2.167e-3 nrs=3.667e-3 sa=440e-9 sb=440e-9
+ sd=520e-9 dtemp=0.0 par=1
C3 n8 DVSS $[nmoscap_6p0] m=8.0 l=10e-6 w=25e-6
R4 n11 n15 $SUB=DVDD $[ppolyf_u] $W=800e-9 $L=63.855e-6 m=1.0 r=29.999e3 par=1
R5 n10 n11 $SUB=DVDD $[ppolyf_u] $W=800e-9 $L=63.855e-6 m=1.0 r=29.999e3 par=1
R6 n19 n10 $SUB=DVDD $[ppolyf_u] $W=800e-9 $L=63.855e-6 m=1.0 r=29.999e3 par=1
R7 n21 n19 $SUB=DVDD $[ppolyf_u] $W=800e-9 $L=63.855e-6 m=1.0 r=29.999e3 par=1
R8 n17 n21 $SUB=DVDD $[ppolyf_u] $W=800e-9 $L=63.855e-6 m=1.0 r=29.999e3 par=1
R9 n20 n8 $SUB=DVDD $[ppolyf_u] $W=800e-9 $L=63.855e-6 m=1.0 r=29.999e3 par=1
R10 n22 n20 $SUB=DVDD $[ppolyf_u] $W=800e-9 $L=63.855e-6 m=1.0 r=29.999e3 par=1
R11 n18 n22 $SUB=DVDD $[ppolyf_u] $W=800e-9 $L=63.855e-6 m=1.0 r=29.999e3 par=1
R12 n13 n18 $SUB=DVDD $[ppolyf_u] $W=800e-9 $L=63.855e-6 m=1.0 r=29.999e3 par=1
R13 n12 n13 $SUB=DVDD $[ppolyf_u] $W=800e-9 $L=63.855e-6 m=1.0 r=29.999e3 par=1
R14 n15 n12 $SUB=DVDD $[ppolyf_u] $W=800e-9 $L=63.855e-6 m=1.0 r=29.999e3 par=1
R15 DVDD n17 $SUB=DVDD $[ppolyf_u] $W=800e-9 $L=63.855e-6 m=1.0 r=29.999e3 par=1
M16 n7 n8 DVSS DVSS nmos_6p0 m=1.0 w=5e-6 l=700e-9 nf=1.0 as=2.2e-12 ad=2.2e-12
+ ps=10.88e-6 pd=10.88e-6 nrd=88e-3 nrs=88e-3 sa=440e-9 sb=440e-9 sd=0.0
+ dtemp=0.0 par=1
M17 DVDD n4 DVSS DVSS nmos_6p0 m=1.0 w=4e-3 l=700e-9 nf=80.0 as=1.058e-9 ad=1.04e-9
+ ps=4.14232e-3 pd=4.0416e-3 nrd=65e-6 nrs=66e-6 sa=440e-9 sb=440e-9 sd=520e-9
+ dtemp=0.0 par=1
M18 n4 n6 DVSS DVSS nmos_6p0 m=1.0 w=30e-6 l=700e-9 nf=1.0 as=13.2e-12 ad=13.2e-12
+ ps=60.88e-6 pd=60.88e-6 nrd=14.667e-3 nrs=14.667e-3 sa=440e-9 sb=440e-9
+ sd=0.0 dtemp=0.0 par=1
M19 n6 n7 DVSS DVSS nmos_6p0 m=1.0 w=30e-6 l=700e-9 nf=1.0 as=13.2e-12 ad=13.2e-12
+ ps=60.88e-6 pd=60.88e-6 nrd=14.667e-3 nrs=14.667e-3 sa=440e-9 sb=440e-9
+ sd=0.0 dtemp=0.0 par=1
D20 DVSS DVDD np_6p0 m=4.0 AREA=40e-12 PJ=82e-6
C21 DVDD DVSS $[nmoscap_6p0] m=4.0 l=15e-6 w=15e-6
.ENDS
