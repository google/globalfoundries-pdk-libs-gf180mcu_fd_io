# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_io__cor
  CLASS ENDCAP BOTTOMLEFT ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_fd_io__cor 0 0 ;
  SIZE 355 BY 355 ;
  SYMMETRY X Y R90 ;
  SITE GF_COR_Site ;
  PIN DVDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal3 ;
        RECT 334 354 341 355 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 354 334 355 341 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 294 354 301 355 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 354 294 355 301 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 278 354 285 355 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 354 278 355 285 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 270 354 277 355 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 354 270 355 277 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 262 354 269 355 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 354 262 355 269 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 214 354 229 355 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 354 214 355 229 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 206 354 213 355 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 354 206 355 213 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 182 354 197 355 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 354 182 355 197 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 166 354 181 355 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 354 166 355 181 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 150 354 165 355 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 354 150 355 165 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 134 354 149 355 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 354 134 355 149 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 118 354 125 355 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 334 354 341 355 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 354 334 355 341 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 294 354 301 355 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 354 294 355 301 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 278 354 285 355 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 354 278 355 285 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 270 354 277 355 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 354 270 355 277 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 262 354 269 355 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 354 262 355 269 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 214 354 229 355 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 354 214 355 229 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 206 354 213 355 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 354 206 355 213 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 182 354 197 355 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 354 182 355 197 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 166 354 181 355 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 354 166 355 181 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 150 354 165 355 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 354 150 355 165 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 134 354 149 355 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 354 134 355 149 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 118 354 125 355 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 354 118 355 125 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 354 118 355 125 ;
    END
  END DVDD
  PIN DVSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal3 ;
        RECT 342 354 348.39 355 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 354 342 355 348.39 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 326 354 333 355 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 354 326 355 333 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 302 354 309 355 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 354 302 355 309 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 286 354 293 355 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 354 286 355 293 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 230 354 245 355 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 354 230 355 245 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 198 354 205 355 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 354 198 355 205 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 126 354 133 355 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 354 126 355 133 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 102 354 117 355 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 354 102 355 117 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 86 354 101 355 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 354 86 355 101 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 70 354 85 355 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 342 354 348.39 355 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 354 342 355 348.39 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 326 354 333 355 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 354 326 355 333 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 302 354 309 355 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 354 302 355 309 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 286 354 293 355 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 354 286 355 293 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 230 354 245 355 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 354 230 355 245 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 198 354 205 355 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 354 198 355 205 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 126 354 133 355 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 354 126 355 133 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 102 354 117 355 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 354 102 355 117 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 86 354 101 355 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 354 86 355 101 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 70 354 85 355 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 354 70 355 85 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 354 70 355 85 ;
    END
  END DVSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal3 ;
        RECT 310 354 317 355 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 354 310 355 317 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 254 354 261 355 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 310 354 317 355 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 354 310 355 317 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 254 354 261 355 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 354 254 355 261 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 354 254 355 261 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal3 ;
        RECT 318 354 325 355 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 354 318 355 325 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 246 354 253 355 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 318 354 325 355 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 354 318 355 325 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 246 354 253 355 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 354 246 355 253 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 354 246 355 253 ;
    END
  END VSS
  OBS
    LAYER Metal1 ;
      RECT 0 0 355 355 ;
    LAYER Metal2 ;
      RECT 0 0 355 355 ;
    LAYER Metal3 ;
      POLYGON 355 69.72 353.72 69.72 353.72 85.28 355 85.28 355 85.72 353.72 85.72 353.72 101.28 355 101.28 355 101.72 353.72 101.72 353.72 117.28 355 117.28 355 117.72 353.72 117.72 353.72 125.28 355 125.28 355 125.72 353.72 125.72 353.72 133.28 355 133.28 355 133.72 353.72 133.72 353.72 149.28 355 149.28 355 149.72 353.72 149.72 353.72 165.28 355 165.28 355 165.72 353.72 165.72 353.72 181.28 355 181.28 355 181.72 353.72 181.72 353.72 197.28 355 197.28 355 197.72 353.72 197.72 353.72 205.28 355 205.28 355 205.72 353.72 205.72 353.72 213.28 355 213.28 355 213.72 353.72 213.72 353.72 229.28 355 229.28 355 229.72 353.72 229.72 353.72 245.28 355 245.28 355 245.72 353.72 245.72 353.72 253.28 355 253.28 355 253.72 353.72 253.72 353.72 261.28 355 261.28 355 261.72 353.72 261.72 353.72 269.28 355 269.28 355 269.72 353.72 269.72 353.72 277.28 355 277.28 355 277.72 353.72 277.72 353.72 285.28 355 285.28 355 285.72 353.72 285.72 353.72 293.28 355 293.28 355 293.72 353.72 293.72 353.72 301.28 355 301.28 355 301.72 353.72 301.72 353.72 309.28 355 309.28 355 309.72 353.72 309.72 353.72 317.28 355 317.28 355 317.72 353.72 317.72 353.72 325.28 355 325.28 355 325.72 353.72 325.72 353.72 333.28 355 333.28 355 333.72 353.72 333.72 353.72 341.28 355 341.28 355 341.72 353.72 341.72 353.72 348.67 355 348.67 355 355 348.67 355 348.67 353.72 341.72 353.72 341.72 355 341.28 355 341.28 353.72 333.72 353.72 333.72 355 333.28 355 333.28 353.72 325.72 353.72 325.72 355 325.28 355 325.28 353.72 317.72 353.72 317.72 355 317.28 355 317.28 353.72 309.72 353.72 309.72 355 309.28 355 309.28 353.72 301.72 353.72 301.72 355 301.28 355 301.28 353.72 293.72 353.72 293.72 355 293.28 355 293.28 353.72 285.72 353.72 285.72 355 285.28 355 285.28 353.72 277.72 353.72 277.72 355 277.28 355 277.28 353.72 269.72 353.72 269.72 355 269.28 355 269.28 353.72 261.72 353.72 261.72 355 261.28 355 261.28 353.72 253.72 353.72 253.72 355 253.28 355 253.28 353.72 245.72 353.72 245.72 355 245.28 355 245.28 353.72 229.72 353.72 229.72 355 229.28 355 229.28 353.72 213.72 353.72 213.72 355 213.28 355 213.28 353.72 205.72 353.72 205.72 355 205.28 355 205.28 353.72 197.72 353.72 197.72 355 197.28 355 197.28 353.72 181.72 353.72 181.72 355 181.28 355 181.28 353.72 165.72 353.72 165.72 355 165.28 355 165.28 353.72 149.72 353.72 149.72 355 149.28 355 149.28 353.72 133.72 353.72 133.72 355 133.28 355 133.28 353.72 125.72 353.72 125.72 355 125.28 355 125.28 353.72 117.72 353.72 117.72 355 117.28 355 117.28 353.72 101.72 353.72 101.72 355 101.28 355 101.28 353.72 85.72 353.72 85.72 355 85.28 355 85.28 353.72 69.72 353.72 69.72 355 0 355 0 0 355 0 ;
    LAYER Metal4 ;
      POLYGON 355 69.72 353.72 69.72 353.72 85.28 355 85.28 355 85.72 353.72 85.72 353.72 101.28 355 101.28 355 101.72 353.72 101.72 353.72 117.28 355 117.28 355 117.72 353.72 117.72 353.72 125.28 355 125.28 355 125.72 353.72 125.72 353.72 133.28 355 133.28 355 133.72 353.72 133.72 353.72 149.28 355 149.28 355 149.72 353.72 149.72 353.72 165.28 355 165.28 355 165.72 353.72 165.72 353.72 181.28 355 181.28 355 181.72 353.72 181.72 353.72 197.28 355 197.28 355 197.72 353.72 197.72 353.72 205.28 355 205.28 355 205.72 353.72 205.72 353.72 213.28 355 213.28 355 213.72 353.72 213.72 353.72 229.28 355 229.28 355 229.72 353.72 229.72 353.72 245.28 355 245.28 355 245.72 353.72 245.72 353.72 253.28 355 253.28 355 253.72 353.72 253.72 353.72 261.28 355 261.28 355 261.72 353.72 261.72 353.72 269.28 355 269.28 355 269.72 353.72 269.72 353.72 277.28 355 277.28 355 277.72 353.72 277.72 353.72 285.28 355 285.28 355 285.72 353.72 285.72 353.72 293.28 355 293.28 355 293.72 353.72 293.72 353.72 301.28 355 301.28 355 301.72 353.72 301.72 353.72 309.28 355 309.28 355 309.72 353.72 309.72 353.72 317.28 355 317.28 355 317.72 353.72 317.72 353.72 325.28 355 325.28 355 325.72 353.72 325.72 353.72 333.28 355 333.28 355 333.72 353.72 333.72 353.72 341.28 355 341.28 355 341.72 353.72 341.72 353.72 348.67 355 348.67 355 355 348.67 355 348.67 353.72 341.72 353.72 341.72 355 341.28 355 341.28 353.72 333.72 353.72 333.72 355 333.28 355 333.28 353.72 325.72 353.72 325.72 355 325.28 355 325.28 353.72 317.72 353.72 317.72 355 317.28 355 317.28 353.72 309.72 353.72 309.72 355 309.28 355 309.28 353.72 301.72 353.72 301.72 355 301.28 355 301.28 353.72 293.72 353.72 293.72 355 293.28 355 293.28 353.72 285.72 353.72 285.72 355 285.28 355 285.28 353.72 277.72 353.72 277.72 355 277.28 355 277.28 353.72 269.72 353.72 269.72 355 269.28 355 269.28 353.72 261.72 353.72 261.72 355 261.28 355 261.28 353.72 253.72 353.72 253.72 355 253.28 355 253.28 353.72 245.72 353.72 245.72 355 245.28 355 245.28 353.72 229.72 353.72 229.72 355 229.28 355 229.28 353.72 213.72 353.72 213.72 355 213.28 355 213.28 353.72 205.72 353.72 205.72 355 205.28 355 205.28 353.72 197.72 353.72 197.72 355 197.28 355 197.28 353.72 181.72 353.72 181.72 355 181.28 355 181.28 353.72 165.72 353.72 165.72 355 165.28 355 165.28 353.72 149.72 353.72 149.72 355 149.28 355 149.28 353.72 133.72 353.72 133.72 355 133.28 355 133.28 353.72 125.72 353.72 125.72 355 125.28 355 125.28 353.72 117.72 353.72 117.72 355 117.28 355 117.28 353.72 101.72 353.72 101.72 355 101.28 355 101.28 353.72 85.72 353.72 85.72 355 85.28 355 85.28 353.72 69.72 353.72 69.72 355 0 355 0 0 355 0 ;
    LAYER Via1 ;
      RECT 0 0 355 355 ;
    LAYER Via2 ;
      RECT 0 0 355 355 ;
    LAYER Via3 ;
      RECT 0 0 355 355 ;
  END

END gf180mcu_fd_io__cor
