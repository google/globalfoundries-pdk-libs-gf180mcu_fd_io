* Copyright 2022 GlobalFoundries PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.SUBCKT gf180mcu_fd_io__in_c DVDD DVSS PAD PD PU VDD VSS Y
C0 DVDD DVSS $[nmoscap_6p0] m=8.0 l=1.5e-6 w=5e-6
C1 DVDD DVSS $[nmoscap_6p0] m=4.0 l=3e-6 w=3e-6
R2 n0 VSS $SUB=VDD $[ppolyf_u] $W=800e-9 $L=3.9e-6 m=1.0 r=1.88247e3 par=1
R3 VDD n6 $SUB=VDD $[ppolyf_u] $W=800e-9 $L=3.9e-6 m=1.0 r=1.88247e3 par=1
M4 n62 n70 DVSS DVSS nmos_6p0 m=1.0 w=3e-6 l=700e-9 nf=1.0 as=1.32e-12 ad=1.32e-12
+ ps=6.88e-6 pd=6.88e-6 nrd=146.667e-3 nrs=146.667e-3 sa=440e-9 sb=440e-9
+ sd=0.0 dtemp=0.0 par=1
M5 n32 n62 DVSS DVSS nmos_6p0 m=1.0 w=3e-6 l=700e-9 nf=1.0 as=1.32e-12 ad=1.32e-12
+ ps=6.88e-6 pd=6.88e-6 nrd=146.667e-3 nrs=146.667e-3 sa=440e-9 sb=440e-9
+ sd=0.0 dtemp=0.0 par=1
M6 n67 n0 VSS VSS nmos_6p0 m=1.0 w=3e-6 l=700e-9 nf=1.0 as=1.32e-12 ad=1.32e-12
+ ps=6.88e-6 pd=6.88e-6 nrd=146.667e-3 nrs=146.667e-3 sa=440e-9 sb=440e-9
+ sd=0.0 dtemp=0.0 par=1
M7 n70 n0 n67 VSS nmos_6p0 m=1.0 w=3e-6 l=700e-9 nf=1.0 as=1.32e-12 ad=1.32e-12
+ ps=6.88e-6 pd=6.88e-6 nrd=146.667e-3 nrs=146.667e-3 sa=440e-9 sb=440e-9
+ sd=0.0 dtemp=0.0 par=1
M8 n62 n70 DVDD DVDD pmos_6p0 m=1.0 w=6e-6 l=700e-9 nf=1.0 as=2.64e-12 ad=2.64e-12
+ ps=12.88e-6 pd=12.88e-6 nrd=73.333e-3 nrs=73.333e-3 sa=440e-9 sb=440e-9
+ sd=0.0 dtemp=0.0 par=1
M9 n32 n62 DVDD DVDD pmos_6p0 m=1.0 w=6e-6 l=700e-9 nf=1.0 as=2.64e-12 ad=2.64e-12
+ ps=12.88e-6 pd=12.88e-6 nrd=73.333e-3 nrs=73.333e-3 sa=440e-9 sb=440e-9
+ sd=0.0 dtemp=0.0 par=1
M10 n70 n0 VDD VDD pmos_6p0 m=1.0 w=3e-6 l=700e-9 nf=1.0 as=1.32e-12 ad=1.32e-12
+ ps=6.88e-6 pd=6.88e-6 nrd=146.667e-3 nrs=146.667e-3 sa=440e-9 sb=440e-9
+ sd=0.0 dtemp=0.0 par=1
M11 n70 n0 VDD VDD pmos_6p0 m=1.0 w=3e-6 l=700e-9 nf=1.0 as=1.32e-12 ad=1.32e-12
+ ps=6.88e-6 pd=6.88e-6 nrd=146.667e-3 nrs=146.667e-3 sa=440e-9 sb=440e-9
+ sd=0.0 dtemp=0.0 par=1
M12 PAD n38 DVDD DVDD pmos_6p0_sab m=1.0 w=80e-6 l=700e-9 nf=2.0 s_sab=280e-9
+ d_sab=2.78e-6 par=1 dtemp=0.0
M13 PAD n50 DVSS DVSS nmos_6p0_sab m=1.0 w=38e-6 l=1.15e-6 nf=1.0 s_sab=280e-9
+ d_sab=3.78e-6 par=1 dtemp=0.0
M14 PAD n47 DVSS DVSS nmos_6p0_sab m=1.0 w=38e-6 l=1.15e-6 nf=1.0 s_sab=280e-9
+ d_sab=3.78e-6 par=1 dtemp=0.0
M15 PAD n43 DVDD DVDD pmos_6p0_sab m=1.0 w=40e-6 l=700e-9 nf=1.0 s_sab=280e-9
+ d_sab=2.78e-6 par=1 dtemp=0.0
M16 PAD n37 DVDD DVDD pmos_6p0_sab m=1.0 w=80e-6 l=700e-9 nf=2.0 s_sab=280e-9
+ d_sab=2.78e-6 par=1 dtemp=0.0
M17 PAD n51 DVSS DVSS nmos_6p0_sab m=1.0 w=38e-6 l=1.15e-6 nf=1.0 s_sab=280e-9
+ d_sab=3.78e-6 par=1 dtemp=0.0
M18 PAD n46 DVSS DVSS nmos_6p0_sab m=1.0 w=38e-6 l=1.15e-6 nf=1.0 s_sab=280e-9
+ d_sab=3.78e-6 par=1 dtemp=0.0
M19 PAD n42 DVDD DVDD pmos_6p0_sab m=1.0 w=40e-6 l=700e-9 nf=1.0 s_sab=280e-9
+ d_sab=2.78e-6 par=1 dtemp=0.0
M20 PAD n39 DVDD DVDD pmos_6p0_sab m=1.0 w=80e-6 l=700e-9 nf=2.0 s_sab=280e-9
+ d_sab=2.78e-6 par=1 dtemp=0.0
M21 PAD n49 DVSS DVSS nmos_6p0_sab m=1.0 w=38e-6 l=1.15e-6 nf=1.0 s_sab=280e-9
+ d_sab=3.78e-6 par=1 dtemp=0.0
M22 PAD n48 DVSS DVSS nmos_6p0_sab m=1.0 w=38e-6 l=1.15e-6 nf=1.0 s_sab=280e-9
+ d_sab=3.78e-6 par=1 dtemp=0.0
M23 PAD n44 DVDD DVDD pmos_6p0_sab m=1.0 w=40e-6 l=700e-9 nf=1.0 s_sab=280e-9
+ d_sab=2.78e-6 par=1 dtemp=0.0
M24 PAD n40 DVDD DVDD pmos_6p0_sab m=1.0 w=80e-6 l=700e-9 nf=2.0 s_sab=280e-9
+ d_sab=2.78e-6 par=1 dtemp=0.0
M25 PAD n52 DVSS DVSS nmos_6p0_sab m=1.0 w=38e-6 l=1.15e-6 nf=1.0 s_sab=280e-9
+ d_sab=3.78e-6 par=1 dtemp=0.0
M26 PAD n45 DVSS DVSS nmos_6p0_sab m=1.0 w=38e-6 l=1.15e-6 nf=1.0 s_sab=280e-9
+ d_sab=3.78e-6 par=1 dtemp=0.0
M27 PAD n41 DVDD DVDD pmos_6p0_sab m=1.0 w=40e-6 l=700e-9 nf=1.0 s_sab=280e-9
+ d_sab=2.78e-6 par=1 dtemp=0.0
M28 n53 n36 DVSS DVSS nmos_6p0 m=1.0 w=3e-6 l=700e-9 nf=2.0 as=1.32e-12 ad=780e-15
+ ps=7.76e-6 pd=4.04e-6 nrd=86.667e-3 nrs=146.667e-3 sa=440e-9 sb=440e-9
+ sd=520e-9 dtemp=0.0 par=1
M29 n170 n0 VSS VSS nmos_6p0 m=1.0 w=1.5e-6 l=700e-9 nf=1.0 as=660e-15
+ ad=660e-15 ps=3.88e-6 pd=3.88e-6 nrd=293.333e-3 nrs=293.333e-3 sa=440e-9
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M30 n36 n170 DVSS DVSS nmos_6p0 m=1.0 w=3e-6 l=700e-9 nf=2.0 as=1.32e-12
+ ad=780e-15 ps=7.76e-6 pd=4.04e-6 nrd=86.667e-3 nrs=146.667e-3 sa=440e-9
+ sb=440e-9 sd=520e-9 dtemp=0.0 par=1
M31 n53 n36 DVDD DVDD pmos_6p0 m=1.0 w=6e-6 l=700e-9 nf=2.0 as=2.64e-12
+ ad=1.56e-12 ps=13.76e-6 pd=7.04e-6 nrd=43.333e-3 nrs=73.333e-3 sa=440e-9
+ sb=440e-9 sd=520e-9 dtemp=0.0 par=1
M32 n170 n0 VDD VDD pmos_6p0 m=1.0 w=3e-6 l=700e-9 nf=1.0 as=1.32e-12
+ ad=1.32e-12 ps=6.88e-6 pd=6.88e-6 nrd=146.667e-3 nrs=146.667e-3 sa=440e-9
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M33 n36 n170 DVDD DVDD pmos_6p0 m=1.0 w=6e-6 l=700e-9 nf=2.0 as=2.64e-12
+ ad=1.56e-12 ps=13.76e-6 pd=7.04e-6 nrd=43.333e-3 nrs=73.333e-3 sa=440e-9
+ sb=440e-9 sd=520e-9 dtemp=0.0 par=1
D34 n0 VDD pn_6p0 m=1.0 AREA=1e-12 PJ=4e-6
D35 n0 VDD pn_6p0 m=1.0 AREA=1e-12 PJ=4e-6
D36 VSS n0 pn_6p0 m=1.0 AREA=230.4e-15 PJ=1.92e-6
D37 VSS n0 pn_6p0 m=1.0 AREA=230.4e-15 PJ=1.92e-6
M38 n183 n0 VSS VSS nmos_6p0 m=1.0 w=3e-6 l=700e-9 nf=1.0 as=1.32e-12
+ ad=1.32e-12 ps=6.88e-6 pd=6.88e-6 nrd=146.667e-3 nrs=146.667e-3 sa=440e-9
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M39 n174 n0 n183 VSS nmos_6p0 m=1.0 w=3e-6 l=700e-9 nf=1.0 as=1.32e-12
+ ad=1.32e-12 ps=6.88e-6 pd=6.88e-6 nrd=146.667e-3 nrs=146.667e-3 sa=440e-9
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M40 n34 n31 DVSS DVSS nmos_6p0 m=1.0 w=3e-6 l=700e-9 nf=1.0 as=1.32e-12
+ ad=1.32e-12 ps=6.88e-6 pd=6.88e-6 nrd=146.667e-3 nrs=146.667e-3 sa=440e-9
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M41 n31 n174 DVSS DVSS nmos_6p0 m=1.0 w=3e-6 l=700e-9 nf=1.0 as=1.32e-12
+ ad=1.32e-12 ps=6.88e-6 pd=6.88e-6 nrd=146.667e-3 nrs=146.667e-3 sa=440e-9
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M42 n174 n0 VDD VDD pmos_6p0 m=1.0 w=3e-6 l=700e-9 nf=1.0 as=1.32e-12
+ ad=1.32e-12 ps=6.88e-6 pd=6.88e-6 nrd=146.667e-3 nrs=146.667e-3 sa=440e-9
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M43 n174 n0 VDD VDD pmos_6p0 m=1.0 w=3e-6 l=700e-9 nf=1.0 as=1.32e-12
+ ad=1.32e-12 ps=6.88e-6 pd=6.88e-6 nrd=146.667e-3 nrs=146.667e-3 sa=440e-9
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M44 n34 n31 DVDD DVDD pmos_6p0 m=1.0 w=6e-6 l=700e-9 nf=1.0 as=2.64e-12
+ ad=2.64e-12 ps=12.88e-6 pd=12.88e-6 nrd=73.333e-3 nrs=73.333e-3 sa=440e-9
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M45 n31 n174 DVDD DVDD pmos_6p0 m=1.0 w=6e-6 l=700e-9 nf=1.0 as=2.64e-12
+ ad=2.64e-12 ps=12.88e-6 pd=12.88e-6 nrd=73.333e-3 nrs=73.333e-3 sa=440e-9
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
D46 VSS n0 pn_6p0 m=1.0 AREA=230.4e-15 PJ=1.92e-6
D47 VSS n0 pn_6p0 m=1.0 AREA=230.4e-15 PJ=1.92e-6
M48 n193 n0 VSS VSS nmos_6p0 m=1.0 w=3e-6 l=700e-9 nf=1.0 as=1.32e-12
+ ad=1.32e-12 ps=6.88e-6 pd=6.88e-6 nrd=146.667e-3 nrs=146.667e-3 sa=440e-9
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M49 n184 n0 n193 VSS nmos_6p0 m=1.0 w=3e-6 l=700e-9 nf=1.0 as=1.32e-12
+ ad=1.32e-12 ps=6.88e-6 pd=6.88e-6 nrd=146.667e-3 nrs=146.667e-3 sa=440e-9
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M50 n30 n28 DVSS DVSS nmos_6p0 m=1.0 w=3e-6 l=700e-9 nf=1.0 as=1.32e-12
+ ad=1.32e-12 ps=6.88e-6 pd=6.88e-6 nrd=146.667e-3 nrs=146.667e-3 sa=440e-9
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M51 n28 n184 DVSS DVSS nmos_6p0 m=1.0 w=3e-6 l=700e-9 nf=1.0 as=1.32e-12
+ ad=1.32e-12 ps=6.88e-6 pd=6.88e-6 nrd=146.667e-3 nrs=146.667e-3 sa=440e-9
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M52 n184 n0 VDD VDD pmos_6p0 m=1.0 w=3e-6 l=700e-9 nf=1.0 as=1.32e-12
+ ad=1.32e-12 ps=6.88e-6 pd=6.88e-6 nrd=146.667e-3 nrs=146.667e-3 sa=440e-9
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M53 n184 n0 VDD VDD pmos_6p0 m=1.0 w=3e-6 l=700e-9 nf=1.0 as=1.32e-12
+ ad=1.32e-12 ps=6.88e-6 pd=6.88e-6 nrd=146.667e-3 nrs=146.667e-3 sa=440e-9
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M54 n30 n28 DVDD DVDD pmos_6p0 m=1.0 w=6e-6 l=700e-9 nf=1.0 as=2.64e-12
+ ad=2.64e-12 ps=12.88e-6 pd=12.88e-6 nrd=73.333e-3 nrs=73.333e-3 sa=440e-9
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M55 n28 n184 DVDD DVDD pmos_6p0 m=1.0 w=6e-6 l=700e-9 nf=1.0 as=2.64e-12
+ ad=2.64e-12 ps=12.88e-6 pd=12.88e-6 nrd=73.333e-3 nrs=73.333e-3 sa=440e-9
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
D56 VSS VDD pn_6p0 m=1.0 AREA=230.4e-15 PJ=1.92e-6
D57 VSS n0 pn_6p0 m=1.0 AREA=230.4e-15 PJ=1.92e-6
M58 n203 VDD VSS VSS nmos_6p0 m=1.0 w=3e-6 l=700e-9 nf=1.0 as=1.32e-12
+ ad=1.32e-12 ps=6.88e-6 pd=6.88e-6 nrd=146.667e-3 nrs=146.667e-3 sa=440e-9
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M59 n194 n0 n203 VSS nmos_6p0 m=1.0 w=3e-6 l=700e-9 nf=1.0 as=1.32e-12
+ ad=1.32e-12 ps=6.88e-6 pd=6.88e-6 nrd=146.667e-3 nrs=146.667e-3 sa=440e-9
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M60 n27 n26 DVSS DVSS nmos_6p0 m=1.0 w=3e-6 l=700e-9 nf=1.0 as=1.32e-12
+ ad=1.32e-12 ps=6.88e-6 pd=6.88e-6 nrd=146.667e-3 nrs=146.667e-3 sa=440e-9
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M61 n26 n194 DVSS DVSS nmos_6p0 m=1.0 w=3e-6 l=700e-9 nf=1.0 as=1.32e-12
+ ad=1.32e-12 ps=6.88e-6 pd=6.88e-6 nrd=146.667e-3 nrs=146.667e-3 sa=440e-9
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M62 n194 VDD VDD VDD pmos_6p0 m=1.0 w=3e-6 l=700e-9 nf=1.0 as=1.32e-12
+ ad=1.32e-12 ps=6.88e-6 pd=6.88e-6 nrd=146.667e-3 nrs=146.667e-3 sa=440e-9
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M63 n194 n0 VDD VDD pmos_6p0 m=1.0 w=3e-6 l=700e-9 nf=1.0 as=1.32e-12
+ ad=1.32e-12 ps=6.88e-6 pd=6.88e-6 nrd=146.667e-3 nrs=146.667e-3 sa=440e-9
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M64 n27 n26 DVDD DVDD pmos_6p0 m=1.0 w=6e-6 l=700e-9 nf=1.0 as=2.64e-12
+ ad=2.64e-12 ps=12.88e-6 pd=12.88e-6 nrd=73.333e-3 nrs=73.333e-3 sa=440e-9
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M65 n26 n194 DVDD DVDD pmos_6p0 m=1.0 w=6e-6 l=700e-9 nf=1.0 as=2.64e-12
+ ad=2.64e-12 ps=12.88e-6 pd=12.88e-6 nrd=73.333e-3 nrs=73.333e-3 sa=440e-9
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M66 n41 n53 n40 DVSS nmos_6p0 m=1.0 w=12e-6 l=700e-9 nf=1.0 as=5.28e-12
+ ad=5.28e-12 ps=24.88e-6 pd=24.88e-6 nrd=36.667e-3 nrs=36.667e-3 sa=440e-9
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M67 n40 DVDD n41 DVSS nmos_6p0 m=1.0 w=1.2e-6 l=700e-9 nf=1.0 as=528e-15
+ ad=528e-15 ps=3.28e-6 pd=3.28e-6 nrd=366.667e-3 nrs=366.667e-3 sa=440e-9
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M68 n45 n204 DVSS DVSS nmos_6p0 m=1.0 w=12e-6 l=700e-9 nf=1.0 as=5.28e-12
+ ad=5.28e-12 ps=24.88e-6 pd=24.88e-6 nrd=36.667e-3 nrs=36.667e-3 sa=440e-9
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M69 n52 n204 DVSS DVSS nmos_6p0 m=1.0 w=12e-6 l=700e-9 nf=1.0 as=5.28e-12
+ ad=5.28e-12 ps=24.88e-6 pd=24.88e-6 nrd=36.667e-3 nrs=36.667e-3 sa=440e-9
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M70 n41 n209 DVSS DVSS nmos_6p0 m=1.0 w=12e-6 l=700e-9 nf=1.0 as=5.28e-12
+ ad=5.28e-12 ps=24.88e-6 pd=24.88e-6 nrd=36.667e-3 nrs=36.667e-3 sa=440e-9
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M71 n209 n32 DVSS DVSS nmos_6p0 m=1.0 w=6e-6 l=700e-9 nf=1.0 as=2.64e-12
+ ad=2.64e-12 ps=12.88e-6 pd=12.88e-6 nrd=73.333e-3 nrs=73.333e-3 sa=440e-9
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M72 n209 n34 DVSS DVSS nmos_6p0 m=1.0 w=6e-6 l=700e-9 nf=1.0 as=2.64e-12
+ ad=2.64e-12 ps=12.88e-6 pd=12.88e-6 nrd=73.333e-3 nrs=73.333e-3 sa=440e-9
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M73 n204 n31 n209 DVSS nmos_6p0 m=1.0 w=6e-6 l=700e-9 nf=1.0 as=2.64e-12
+ ad=2.64e-12 ps=12.88e-6 pd=12.88e-6 nrd=73.333e-3 nrs=73.333e-3 sa=440e-9
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M74 n45 n36 n52 DVDD pmos_6p0 m=1.0 w=24e-6 l=700e-9 nf=1.0 as=10.56e-12
+ ad=10.56e-12 ps=48.88e-6 pd=48.88e-6 nrd=18.333e-3 nrs=18.333e-3 sa=440e-9
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M75 n204 n31 DVDD DVDD pmos_6p0 m=1.0 w=12e-6 l=700e-9 nf=1.0 as=5.28e-12
+ ad=5.28e-12 ps=24.88e-6 pd=24.88e-6 nrd=36.667e-3 nrs=36.667e-3 sa=440e-9
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M76 n41 n209 DVDD DVDD pmos_6p0 m=1.0 w=24e-6 l=700e-9 nf=1.0 as=10.56e-12
+ ad=10.56e-12 ps=48.88e-6 pd=48.88e-6 nrd=18.333e-3 nrs=18.333e-3 sa=440e-9
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M77 n52 n204 DVDD DVDD pmos_6p0 m=1.0 w=24e-6 l=700e-9 nf=1.0 as=10.56e-12
+ ad=10.56e-12 ps=48.88e-6 pd=48.88e-6 nrd=18.333e-3 nrs=18.333e-3 sa=440e-9
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M78 n45 DVSS n52 DVDD pmos_6p0 m=1.0 w=1.2e-6 l=700e-9 nf=1.0 as=528e-15
+ ad=528e-15 ps=3.28e-6 pd=3.28e-6 nrd=366.667e-3 nrs=366.667e-3 sa=440e-9
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M79 n204 n32 DVDD DVDD pmos_6p0 m=1.0 w=12e-6 l=700e-9 nf=1.0 as=5.28e-12
+ ad=5.28e-12 ps=24.88e-6 pd=24.88e-6 nrd=36.667e-3 nrs=36.667e-3 sa=440e-9
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M80 n209 n34 n204 DVDD pmos_6p0 m=1.0 w=12e-6 l=700e-9 nf=1.0 as=5.28e-12
+ ad=5.28e-12 ps=24.88e-6 pd=24.88e-6 nrd=36.667e-3 nrs=36.667e-3 sa=440e-9
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M81 n40 n209 DVDD DVDD pmos_6p0 m=1.0 w=24e-6 l=700e-9 nf=1.0 as=10.56e-12
+ ad=10.56e-12 ps=48.88e-6 pd=48.88e-6 nrd=18.333e-3 nrs=18.333e-3 sa=440e-9
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M82 n42 n53 n37 DVSS nmos_6p0 m=1.0 w=12e-6 l=700e-9 nf=1.0 as=5.28e-12
+ ad=5.28e-12 ps=24.88e-6 pd=24.88e-6 nrd=36.667e-3 nrs=36.667e-3 sa=440e-9
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M83 n37 DVDD n42 DVSS nmos_6p0 m=1.0 w=1.2e-6 l=700e-9 nf=1.0 as=528e-15
+ ad=528e-15 ps=3.28e-6 pd=3.28e-6 nrd=366.667e-3 nrs=366.667e-3 sa=440e-9
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M84 n46 n217 DVSS DVSS nmos_6p0 m=1.0 w=12e-6 l=700e-9 nf=1.0 as=5.28e-12
+ ad=5.28e-12 ps=24.88e-6 pd=24.88e-6 nrd=36.667e-3 nrs=36.667e-3 sa=440e-9
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M85 n51 n217 DVSS DVSS nmos_6p0 m=1.0 w=12e-6 l=700e-9 nf=1.0 as=5.28e-12
+ ad=5.28e-12 ps=24.88e-6 pd=24.88e-6 nrd=36.667e-3 nrs=36.667e-3 sa=440e-9
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M86 n42 n222 DVSS DVSS nmos_6p0 m=1.0 w=12e-6 l=700e-9 nf=1.0 as=5.28e-12
+ ad=5.28e-12 ps=24.88e-6 pd=24.88e-6 nrd=36.667e-3 nrs=36.667e-3 sa=440e-9
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M87 n222 n32 DVSS DVSS nmos_6p0 m=1.0 w=6e-6 l=700e-9 nf=1.0 as=2.64e-12
+ ad=2.64e-12 ps=12.88e-6 pd=12.88e-6 nrd=73.333e-3 nrs=73.333e-3 sa=440e-9
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M88 n222 n30 DVSS DVSS nmos_6p0 m=1.0 w=6e-6 l=700e-9 nf=1.0 as=2.64e-12
+ ad=2.64e-12 ps=12.88e-6 pd=12.88e-6 nrd=73.333e-3 nrs=73.333e-3 sa=440e-9
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M89 n217 n28 n222 DVSS nmos_6p0 m=1.0 w=6e-6 l=700e-9 nf=1.0 as=2.64e-12
+ ad=2.64e-12 ps=12.88e-6 pd=12.88e-6 nrd=73.333e-3 nrs=73.333e-3 sa=440e-9
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M90 n46 n36 n51 DVDD pmos_6p0 m=1.0 w=24e-6 l=700e-9 nf=1.0 as=10.56e-12
+ ad=10.56e-12 ps=48.88e-6 pd=48.88e-6 nrd=18.333e-3 nrs=18.333e-3 sa=440e-9
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M91 n217 n28 DVDD DVDD pmos_6p0 m=1.0 w=12e-6 l=700e-9 nf=1.0 as=5.28e-12
+ ad=5.28e-12 ps=24.88e-6 pd=24.88e-6 nrd=36.667e-3 nrs=36.667e-3 sa=440e-9
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M92 n42 n222 DVDD DVDD pmos_6p0 m=1.0 w=24e-6 l=700e-9 nf=1.0 as=10.56e-12
+ ad=10.56e-12 ps=48.88e-6 pd=48.88e-6 nrd=18.333e-3 nrs=18.333e-3 sa=440e-9
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M93 n51 n217 DVDD DVDD pmos_6p0 m=1.0 w=24e-6 l=700e-9 nf=1.0 as=10.56e-12
+ ad=10.56e-12 ps=48.88e-6 pd=48.88e-6 nrd=18.333e-3 nrs=18.333e-3 sa=440e-9
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M94 n46 DVSS n51 DVDD pmos_6p0 m=1.0 w=1.2e-6 l=700e-9 nf=1.0 as=528e-15
+ ad=528e-15 ps=3.28e-6 pd=3.28e-6 nrd=366.667e-3 nrs=366.667e-3 sa=440e-9
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M95 n217 n32 DVDD DVDD pmos_6p0 m=1.0 w=12e-6 l=700e-9 nf=1.0 as=5.28e-12
+ ad=5.28e-12 ps=24.88e-6 pd=24.88e-6 nrd=36.667e-3 nrs=36.667e-3 sa=440e-9
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M96 n222 n30 n217 DVDD pmos_6p0 m=1.0 w=12e-6 l=700e-9 nf=1.0 as=5.28e-12
+ ad=5.28e-12 ps=24.88e-6 pd=24.88e-6 nrd=36.667e-3 nrs=36.667e-3 sa=440e-9
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M97 n37 n222 DVDD DVDD pmos_6p0 m=1.0 w=24e-6 l=700e-9 nf=1.0 as=10.56e-12
+ ad=10.56e-12 ps=48.88e-6 pd=48.88e-6 nrd=18.333e-3 nrs=18.333e-3 sa=440e-9
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M98 n43 n53 n38 DVSS nmos_6p0 m=1.0 w=12e-6 l=700e-9 nf=1.0 as=5.28e-12
+ ad=5.28e-12 ps=24.88e-6 pd=24.88e-6 nrd=36.667e-3 nrs=36.667e-3 sa=440e-9
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M99 n38 DVDD n43 DVSS nmos_6p0 m=1.0 w=1.2e-6 l=700e-9 nf=1.0 as=528e-15
+ ad=528e-15 ps=3.28e-6 pd=3.28e-6 nrd=366.667e-3 nrs=366.667e-3 sa=440e-9
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M100 n47 n230 DVSS DVSS nmos_6p0 m=1.0 w=12e-6 l=700e-9 nf=1.0 as=5.28e-12
+ ad=5.28e-12 ps=24.88e-6 pd=24.88e-6 nrd=36.667e-3 nrs=36.667e-3 sa=440e-9
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M101 n50 n230 DVSS DVSS nmos_6p0 m=1.0 w=12e-6 l=700e-9 nf=1.0 as=5.28e-12
+ ad=5.28e-12 ps=24.88e-6 pd=24.88e-6 nrd=36.667e-3 nrs=36.667e-3 sa=440e-9
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M102 n43 n235 DVSS DVSS nmos_6p0 m=1.0 w=12e-6 l=700e-9 nf=1.0 as=5.28e-12
+ ad=5.28e-12 ps=24.88e-6 pd=24.88e-6 nrd=36.667e-3 nrs=36.667e-3 sa=440e-9
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M103 n235 n32 DVSS DVSS nmos_6p0 m=1.0 w=6e-6 l=700e-9 nf=1.0 as=2.64e-12
+ ad=2.64e-12 ps=12.88e-6 pd=12.88e-6 nrd=73.333e-3 nrs=73.333e-3 sa=440e-9
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M104 n235 n30 DVSS DVSS nmos_6p0 m=1.0 w=6e-6 l=700e-9 nf=1.0 as=2.64e-12
+ ad=2.64e-12 ps=12.88e-6 pd=12.88e-6 nrd=73.333e-3 nrs=73.333e-3 sa=440e-9
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M105 n230 n28 n235 DVSS nmos_6p0 m=1.0 w=6e-6 l=700e-9 nf=1.0 as=2.64e-12
+ ad=2.64e-12 ps=12.88e-6 pd=12.88e-6 nrd=73.333e-3 nrs=73.333e-3 sa=440e-9
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M106 n47 n36 n50 DVDD pmos_6p0 m=1.0 w=24e-6 l=700e-9 nf=1.0 as=10.56e-12
+ ad=10.56e-12 ps=48.88e-6 pd=48.88e-6 nrd=18.333e-3 nrs=18.333e-3 sa=440e-9
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M107 n230 n28 DVDD DVDD pmos_6p0 m=1.0 w=12e-6 l=700e-9 nf=1.0 as=5.28e-12
+ ad=5.28e-12 ps=24.88e-6 pd=24.88e-6 nrd=36.667e-3 nrs=36.667e-3 sa=440e-9
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M108 n43 n235 DVDD DVDD pmos_6p0 m=1.0 w=24e-6 l=700e-9 nf=1.0 as=10.56e-12
+ ad=10.56e-12 ps=48.88e-6 pd=48.88e-6 nrd=18.333e-3 nrs=18.333e-3 sa=440e-9
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M109 n50 n230 DVDD DVDD pmos_6p0 m=1.0 w=24e-6 l=700e-9 nf=1.0 as=10.56e-12
+ ad=10.56e-12 ps=48.88e-6 pd=48.88e-6 nrd=18.333e-3 nrs=18.333e-3 sa=440e-9
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M110 n47 DVSS n50 DVDD pmos_6p0 m=1.0 w=1.2e-6 l=700e-9 nf=1.0 as=528e-15
+ ad=528e-15 ps=3.28e-6 pd=3.28e-6 nrd=366.667e-3 nrs=366.667e-3 sa=440e-9
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M111 n230 n32 DVDD DVDD pmos_6p0 m=1.0 w=12e-6 l=700e-9 nf=1.0 as=5.28e-12
+ ad=5.28e-12 ps=24.88e-6 pd=24.88e-6 nrd=36.667e-3 nrs=36.667e-3 sa=440e-9
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M112 n235 n30 n230 DVDD pmos_6p0 m=1.0 w=12e-6 l=700e-9 nf=1.0 as=5.28e-12
+ ad=5.28e-12 ps=24.88e-6 pd=24.88e-6 nrd=36.667e-3 nrs=36.667e-3 sa=440e-9
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M113 n38 n235 DVDD DVDD pmos_6p0 m=1.0 w=24e-6 l=700e-9 nf=1.0 as=10.56e-12
+ ad=10.56e-12 ps=48.88e-6 pd=48.88e-6 nrd=18.333e-3 nrs=18.333e-3 sa=440e-9
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M114 n44 n53 n39 DVSS nmos_6p0 m=1.0 w=12e-6 l=700e-9 nf=1.0 as=5.28e-12
+ ad=5.28e-12 ps=24.88e-6 pd=24.88e-6 nrd=36.667e-3 nrs=36.667e-3 sa=440e-9
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M115 n39 DVDD n44 DVSS nmos_6p0 m=1.0 w=1.2e-6 l=700e-9 nf=1.0 as=528e-15
+ ad=528e-15 ps=3.28e-6 pd=3.28e-6 nrd=366.667e-3 nrs=366.667e-3 sa=440e-9
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M116 n48 n243 DVSS DVSS nmos_6p0 m=1.0 w=12e-6 l=700e-9 nf=1.0 as=5.28e-12
+ ad=5.28e-12 ps=24.88e-6 pd=24.88e-6 nrd=36.667e-3 nrs=36.667e-3 sa=440e-9
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M117 n49 n243 DVSS DVSS nmos_6p0 m=1.0 w=12e-6 l=700e-9 nf=1.0 as=5.28e-12
+ ad=5.28e-12 ps=24.88e-6 pd=24.88e-6 nrd=36.667e-3 nrs=36.667e-3 sa=440e-9
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M118 n44 n248 DVSS DVSS nmos_6p0 m=1.0 w=12e-6 l=700e-9 nf=1.0 as=5.28e-12
+ ad=5.28e-12 ps=24.88e-6 pd=24.88e-6 nrd=36.667e-3 nrs=36.667e-3 sa=440e-9
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M119 n248 n32 DVSS DVSS nmos_6p0 m=1.0 w=6e-6 l=700e-9 nf=1.0 as=2.64e-12
+ ad=2.64e-12 ps=12.88e-6 pd=12.88e-6 nrd=73.333e-3 nrs=73.333e-3 sa=440e-9
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M120 n248 n27 DVSS DVSS nmos_6p0 m=1.0 w=6e-6 l=700e-9 nf=1.0 as=2.64e-12
+ ad=2.64e-12 ps=12.88e-6 pd=12.88e-6 nrd=73.333e-3 nrs=73.333e-3 sa=440e-9
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M121 n243 n26 n248 DVSS nmos_6p0 m=1.0 w=6e-6 l=700e-9 nf=1.0 as=2.64e-12
+ ad=2.64e-12 ps=12.88e-6 pd=12.88e-6 nrd=73.333e-3 nrs=73.333e-3 sa=440e-9
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M122 n48 n36 n49 DVDD pmos_6p0 m=1.0 w=24e-6 l=700e-9 nf=1.0 as=10.56e-12
+ ad=10.56e-12 ps=48.88e-6 pd=48.88e-6 nrd=18.333e-3 nrs=18.333e-3 sa=440e-9
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M123 n243 n26 DVDD DVDD pmos_6p0 m=1.0 w=12e-6 l=700e-9 nf=1.0 as=5.28e-12
+ ad=5.28e-12 ps=24.88e-6 pd=24.88e-6 nrd=36.667e-3 nrs=36.667e-3 sa=440e-9
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M124 n44 n248 DVDD DVDD pmos_6p0 m=1.0 w=24e-6 l=700e-9 nf=1.0 as=10.56e-12
+ ad=10.56e-12 ps=48.88e-6 pd=48.88e-6 nrd=18.333e-3 nrs=18.333e-3 sa=440e-9
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M125 n49 n243 DVDD DVDD pmos_6p0 m=1.0 w=24e-6 l=700e-9 nf=1.0 as=10.56e-12
+ ad=10.56e-12 ps=48.88e-6 pd=48.88e-6 nrd=18.333e-3 nrs=18.333e-3 sa=440e-9
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M126 n48 DVSS n49 DVDD pmos_6p0 m=1.0 w=1.2e-6 l=700e-9 nf=1.0 as=528e-15
+ ad=528e-15 ps=3.28e-6 pd=3.28e-6 nrd=366.667e-3 nrs=366.667e-3 sa=440e-9
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M127 n243 n32 DVDD DVDD pmos_6p0 m=1.0 w=12e-6 l=700e-9 nf=1.0 as=5.28e-12
+ ad=5.28e-12 ps=24.88e-6 pd=24.88e-6 nrd=36.667e-3 nrs=36.667e-3 sa=440e-9
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M128 n248 n27 n243 DVDD pmos_6p0 m=1.0 w=12e-6 l=700e-9 nf=1.0 as=5.28e-12
+ ad=5.28e-12 ps=24.88e-6 pd=24.88e-6 nrd=36.667e-3 nrs=36.667e-3 sa=440e-9
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M129 n39 n248 DVDD DVDD pmos_6p0 m=1.0 w=24e-6 l=700e-9 nf=1.0 as=10.56e-12
+ ad=10.56e-12 ps=48.88e-6 pd=48.88e-6 nrd=18.333e-3 nrs=18.333e-3 sa=440e-9
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M130 n268 n257 DVSS DVSS nmos_6p0 m=1.0 w=3e-6 l=700e-9 nf=2.0 as=1.32e-12
+ ad=780e-15 ps=7.76e-6 pd=4.04e-6 nrd=86.667e-3 nrs=146.667e-3 sa=440e-9
+ sb=440e-9 sd=520e-9 dtemp=0.0 par=1
M131 n281 n6 VSS VSS nmos_6p0 m=1.0 w=1.5e-6 l=700e-9 nf=1.0 as=660e-15
+ ad=660e-15 ps=3.88e-6 pd=3.88e-6 nrd=293.333e-3 nrs=293.333e-3 sa=440e-9
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M132 n257 n281 DVSS DVSS nmos_6p0 m=1.0 w=3e-6 l=700e-9 nf=2.0 as=1.32e-12
+ ad=780e-15 ps=7.76e-6 pd=4.04e-6 nrd=86.667e-3 nrs=146.667e-3 sa=440e-9
+ sb=440e-9 sd=520e-9 dtemp=0.0 par=1
M133 n268 n257 DVDD DVDD pmos_6p0 m=1.0 w=6e-6 l=700e-9 nf=2.0 as=2.64e-12
+ ad=1.56e-12 ps=13.76e-6 pd=7.04e-6 nrd=43.333e-3 nrs=73.333e-3 sa=440e-9
+ sb=440e-9 sd=520e-9 dtemp=0.0 par=1
M134 n281 n6 VDD VDD pmos_6p0 m=1.0 w=3e-6 l=700e-9 nf=1.0 as=1.32e-12
+ ad=1.32e-12 ps=6.88e-6 pd=6.88e-6 nrd=146.667e-3 nrs=146.667e-3 sa=440e-9
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M135 n257 n281 DVDD DVDD pmos_6p0 m=1.0 w=6e-6 l=700e-9 nf=2.0 as=2.64e-12
+ ad=1.56e-12 ps=13.76e-6 pd=7.04e-6 nrd=43.333e-3 nrs=73.333e-3 sa=440e-9
+ sb=440e-9 sd=520e-9 dtemp=0.0 par=1
M136 n274 n258 DVSS DVSS nmos_6p0 m=1.0 w=3e-6 l=700e-9 nf=2.0 as=1.32e-12
+ ad=780e-15 ps=7.76e-6 pd=4.04e-6 nrd=86.667e-3 nrs=146.667e-3 sa=440e-9
+ sb=440e-9 sd=520e-9 dtemp=0.0 par=1
M137 n289 n0 VSS VSS nmos_6p0 m=1.0 w=1.5e-6 l=700e-9 nf=1.0 as=660e-15
+ ad=660e-15 ps=3.88e-6 pd=3.88e-6 nrd=293.333e-3 nrs=293.333e-3 sa=440e-9
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M138 n258 n289 DVSS DVSS nmos_6p0 m=1.0 w=3e-6 l=700e-9 nf=2.0 as=1.32e-12
+ ad=780e-15 ps=7.76e-6 pd=4.04e-6 nrd=86.667e-3 nrs=146.667e-3 sa=440e-9
+ sb=440e-9 sd=520e-9 dtemp=0.0 par=1
M139 n274 n258 DVDD DVDD pmos_6p0 m=1.0 w=6e-6 l=700e-9 nf=2.0 as=2.64e-12
+ ad=1.56e-12 ps=13.76e-6 pd=7.04e-6 nrd=43.333e-3 nrs=73.333e-3 sa=440e-9
+ sb=440e-9 sd=520e-9 dtemp=0.0 par=1
M140 n289 n0 VDD VDD pmos_6p0 m=1.0 w=3e-6 l=700e-9 nf=1.0 as=1.32e-12
+ ad=1.32e-12 ps=6.88e-6 pd=6.88e-6 nrd=146.667e-3 nrs=146.667e-3 sa=440e-9
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M141 n258 n289 DVDD DVDD pmos_6p0 m=1.0 w=6e-6 l=700e-9 nf=2.0 as=2.64e-12
+ ad=1.56e-12 ps=13.76e-6 pd=7.04e-6 nrd=43.333e-3 nrs=73.333e-3 sa=440e-9
+ sb=440e-9 sd=520e-9 dtemp=0.0 par=1
M142 n272 n260 DVSS DVSS nmos_6p0 m=1.0 w=3e-6 l=700e-9 nf=2.0 as=1.32e-12
+ ad=780e-15 ps=7.76e-6 pd=4.04e-6 nrd=86.667e-3 nrs=146.667e-3 sa=440e-9
+ sb=440e-9 sd=520e-9 dtemp=0.0 par=1
M143 n297 n261 VSS VSS nmos_6p0 m=1.0 w=1.5e-6 l=700e-9 nf=1.0 as=660e-15
+ ad=660e-15 ps=3.88e-6 pd=3.88e-6 nrd=293.333e-3 nrs=293.333e-3 sa=440e-9
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M144 n260 n297 DVSS DVSS nmos_6p0 m=1.0 w=3e-6 l=700e-9 nf=2.0 as=1.32e-12
+ ad=780e-15 ps=7.76e-6 pd=4.04e-6 nrd=86.667e-3 nrs=146.667e-3 sa=440e-9
+ sb=440e-9 sd=520e-9 dtemp=0.0 par=1
M145 n272 n260 DVDD DVDD pmos_6p0 m=1.0 w=6e-6 l=700e-9 nf=2.0 as=2.64e-12
+ ad=1.56e-12 ps=13.76e-6 pd=7.04e-6 nrd=43.333e-3 nrs=73.333e-3 sa=440e-9
+ sb=440e-9 sd=520e-9 dtemp=0.0 par=1
M146 n297 n261 VDD VDD pmos_6p0 m=1.0 w=3e-6 l=700e-9 nf=1.0 as=1.32e-12
+ ad=1.32e-12 ps=6.88e-6 pd=6.88e-6 nrd=146.667e-3 nrs=146.667e-3 sa=440e-9
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M147 n260 n297 DVDD DVDD pmos_6p0 m=1.0 w=6e-6 l=700e-9 nf=2.0 as=2.64e-12
+ ad=1.56e-12 ps=13.76e-6 pd=7.04e-6 nrd=43.333e-3 nrs=73.333e-3 sa=440e-9
+ sb=440e-9 sd=520e-9 dtemp=0.0 par=1
M148 n276 n263 DVSS DVSS nmos_6p0 m=1.0 w=3e-6 l=700e-9 nf=2.0 as=1.32e-12
+ ad=780e-15 ps=7.76e-6 pd=4.04e-6 nrd=86.667e-3 nrs=146.667e-3 sa=440e-9
+ sb=440e-9 sd=520e-9 dtemp=0.0 par=1
M149 n305 n259 VSS VSS nmos_6p0 m=1.0 w=1.5e-6 l=700e-9 nf=1.0 as=660e-15
+ ad=660e-15 ps=3.88e-6 pd=3.88e-6 nrd=293.333e-3 nrs=293.333e-3 sa=440e-9
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M150 n263 n305 DVSS DVSS nmos_6p0 m=1.0 w=3e-6 l=700e-9 nf=2.0 as=1.32e-12
+ ad=780e-15 ps=7.76e-6 pd=4.04e-6 nrd=86.667e-3 nrs=146.667e-3 sa=440e-9
+ sb=440e-9 sd=520e-9 dtemp=0.0 par=1
M151 n276 n263 DVDD DVDD pmos_6p0 m=1.0 w=6e-6 l=700e-9 nf=2.0 as=2.64e-12
+ ad=1.56e-12 ps=13.76e-6 pd=7.04e-6 nrd=43.333e-3 nrs=73.333e-3 sa=440e-9
+ sb=440e-9 sd=520e-9 dtemp=0.0 par=1
M152 n305 n259 VDD VDD pmos_6p0 m=1.0 w=3e-6 l=700e-9 nf=1.0 as=1.32e-12
+ ad=1.32e-12 ps=6.88e-6 pd=6.88e-6 nrd=146.667e-3 nrs=146.667e-3 sa=440e-9
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M153 n263 n305 DVDD DVDD pmos_6p0 m=1.0 w=6e-6 l=700e-9 nf=2.0 as=2.64e-12
+ ad=1.56e-12 ps=13.76e-6 pd=7.04e-6 nrd=43.333e-3 nrs=73.333e-3 sa=440e-9
+ sb=440e-9 sd=520e-9 dtemp=0.0 par=1
D154 PD VDD pn_6p0 m=1.0 AREA=1e-12 PJ=4e-6
D155 n6 VDD pn_6p0 m=1.0 AREA=1e-12 PJ=4e-6
D156 n0 VDD pn_6p0 m=1.0 AREA=1e-12 PJ=4e-6
D157 PU VDD pn_6p0 m=1.0 AREA=1e-12 PJ=4e-6
M158 n313 n258 DVDD DVDD pmos_6p0 m=1.0 w=8e-6 l=700e-9 nf=1.0 as=3.52e-12
+ ad=3.52e-12 ps=16.88e-6 pd=16.88e-6 nrd=55e-3 nrs=55e-3 sa=440e-9 sb=440e-9
+ sd=0.0 dtemp=0.0 par=1
M159 DVDD n258 n314 DVDD pmos_6p0 m=1.0 w=3e-6 l=700e-9 nf=1.0 as=1.32e-12
+ ad=1.32e-12 ps=6.88e-6 pd=6.88e-6 nrd=146.667e-3 nrs=146.667e-3 sa=440e-9
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M160 n315 n15 DVDD DVDD pmos_6p0 m=1.0 w=3.8e-6 l=700e-9 nf=1.0 as=1.672e-12
+ ad=1.672e-12 ps=8.48e-6 pd=8.48e-6 nrd=115.789e-3 nrs=115.789e-3 sa=440e-9
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M161 DVSS n314 n315 DVDD pmos_6p0 m=1.0 w=3.8e-6 l=700e-9 nf=1.0 as=1.672e-12
+ ad=1.672e-12 ps=8.48e-6 pd=8.48e-6 nrd=115.789e-3 nrs=115.789e-3 sa=440e-9
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M162 n275 n257 DVDD DVDD pmos_6p0 m=1.0 w=6e-6 l=700e-9 nf=1.0 as=2.64e-12
+ ad=2.64e-12 ps=12.88e-6 pd=12.88e-6 nrd=73.333e-3 nrs=73.333e-3 sa=440e-9
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M163 n275 n313 n310 DVDD pmos_6p0 m=1.0 w=2e-6 l=700e-9 nf=1.0 as=880e-15
+ ad=880e-15 ps=4.88e-6 pd=4.88e-6 nrd=220e-3 nrs=220e-3 sa=440e-9 sb=440e-9
+ sd=0.0 dtemp=0.0 par=1
M164 n275 n313 n314 DVDD pmos_6p0 m=1.0 w=2e-6 l=700e-9 nf=1.0 as=880e-15
+ ad=880e-15 ps=4.88e-6 pd=4.88e-6 nrd=220e-3 nrs=220e-3 sa=440e-9 sb=440e-9
+ sd=0.0 dtemp=0.0 par=1
M165 n275 n15 n315 DVDD pmos_6p0 m=1.0 w=4.3e-6 l=700e-9 nf=1.0 as=1.892e-12
+ ad=1.892e-12 ps=9.48e-6 pd=9.48e-6 nrd=102.326e-3 nrs=102.326e-3 sa=440e-9
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M166 n320 n257 DVSS DVSS nmos_6p0 m=1.0 w=16e-6 l=700e-9 nf=1.0 as=7.04e-12
+ ad=7.04e-12 ps=32.88e-6 pd=32.88e-6 nrd=27.5e-3 nrs=27.5e-3 sa=440e-9
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M167 n312 n15 n320 DVSS nmos_6p0 m=1.0 w=10.6e-6 l=700e-9 nf=1.0 as=4.664e-12
+ ad=4.664e-12 ps=22.08e-6 pd=22.08e-6 nrd=41.509e-3 nrs=41.509e-3 sa=440e-9
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M168 n275 n15 n312 DVSS nmos_6p0 m=1.0 w=12e-6 l=700e-9 nf=1.0 as=5.28e-12
+ ad=5.28e-12 ps=24.88e-6 pd=24.88e-6 nrd=36.667e-3 nrs=36.667e-3 sa=440e-9
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M169 n313 n258 DVSS DVSS nmos_6p0 m=1.0 w=4e-6 l=700e-9 nf=1.0 as=1.76e-12
+ ad=1.76e-12 ps=8.88e-6 pd=8.88e-6 nrd=110e-3 nrs=110e-3 sa=440e-9 sb=440e-9
+ sd=0.0 dtemp=0.0 par=1
M170 n275 n258 n310 DVSS nmos_6p0 m=1.0 w=1.5e-6 l=700e-9 nf=1.0 as=660e-15
+ ad=660e-15 ps=3.88e-6 pd=3.88e-6 nrd=293.333e-3 nrs=293.333e-3 sa=440e-9
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M171 n275 n258 n314 DVSS nmos_6p0 m=1.0 w=1.5e-6 l=700e-9 nf=1.0 as=660e-15
+ ad=660e-15 ps=3.88e-6 pd=3.88e-6 nrd=293.333e-3 nrs=293.333e-3 sa=440e-9
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M172 DVDD n310 n312 DVSS nmos_6p0 m=1.0 w=1.3e-6 l=700e-9 nf=1.0 as=572e-15
+ ad=572e-15 ps=3.48e-6 pd=3.48e-6 nrd=338.462e-3 nrs=338.462e-3 sa=440e-9
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M173 DVSS n313 n310 DVSS nmos_6p0 m=1.0 w=1.5e-6 l=700e-9 nf=1.0 as=660e-15
+ ad=660e-15 ps=3.88e-6 pd=3.88e-6 nrd=293.333e-3 nrs=293.333e-3 sa=440e-9
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M174 n328 n275 DVDD DVDD pmos_6p0 m=1.0 w=2e-6 l=700e-9 nf=1.0 as=880e-15
+ ad=880e-15 ps=4.88e-6 pd=4.88e-6 nrd=220e-3 nrs=220e-3 sa=440e-9 sb=440e-9
+ sd=0.0 dtemp=0.0 par=1
M175 n325 n328 VDD VDD pmos_6p0 m=1.0 w=10e-6 l=700e-9 nf=1.0 as=4.4e-12
+ ad=4.4e-12 ps=20.88e-6 pd=20.88e-6 nrd=44e-3 nrs=44e-3 sa=440e-9 sb=440e-9
+ sd=0.0 dtemp=0.0 par=1
M176 Y n325 VDD VDD pmos_6p0 m=1.0 w=21e-6 l=700e-9 nf=1.0 as=9.24e-12
+ ad=9.24e-12 ps=42.88e-6 pd=42.88e-6 nrd=20.952e-3 nrs=20.952e-3 sa=440e-9
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M177 n328 n275 DVSS DVSS nmos_6p0 m=1.0 w=8e-6 l=700e-9 nf=1.0 as=3.52e-12
+ ad=3.52e-12 ps=16.88e-6 pd=16.88e-6 nrd=55e-3 nrs=55e-3 sa=440e-9 sb=440e-9
+ sd=0.0 dtemp=0.0 par=1
M178 Y n325 VSS VSS nmos_6p0 m=1.0 w=9e-6 l=700e-9 nf=1.0 as=3.96e-12
+ ad=3.96e-12 ps=18.88e-6 pd=18.88e-6 nrd=48.889e-3 nrs=48.889e-3 sa=440e-9
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M179 n325 n328 VSS VSS nmos_6p0 m=1.0 w=2.5e-6 l=700e-9 nf=1.0 as=1.1e-12
+ ad=1.1e-12 ps=5.88e-6 pd=5.88e-6 nrd=176e-3 nrs=176e-3 sa=440e-9 sb=440e-9
+ sd=0.0 dtemp=0.0 par=1
M180 n261 n335 VDD VDD pmos_6p0 m=1.0 w=3e-6 l=700e-9 nf=1.0 as=1.32e-12
+ ad=1.32e-12 ps=6.88e-6 pd=6.88e-6 nrd=146.667e-3 nrs=146.667e-3 sa=440e-9
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M181 n261 PU VDD VDD pmos_6p0 m=1.0 w=3e-6 l=700e-9 nf=1.0 as=1.32e-12
+ ad=1.32e-12 ps=6.88e-6 pd=6.88e-6 nrd=146.667e-3 nrs=146.667e-3 sa=440e-9
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M182 n336 PU VSS VSS nmos_6p0 m=1.0 w=3e-6 l=700e-9 nf=1.0 as=1.32e-12
+ ad=1.32e-12 ps=6.88e-6 pd=6.88e-6 nrd=146.667e-3 nrs=146.667e-3 sa=440e-9
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M183 n261 n335 n336 VSS nmos_6p0 m=1.0 w=3e-6 l=700e-9 nf=1.0 as=1.32e-12
+ ad=1.32e-12 ps=6.88e-6 pd=6.88e-6 nrd=146.667e-3 nrs=146.667e-3 sa=440e-9
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M184 n259 PD VDD VDD pmos_6p0 m=1.0 w=3e-6 l=700e-9 nf=1.0 as=1.32e-12
+ ad=1.32e-12 ps=6.88e-6 pd=6.88e-6 nrd=146.667e-3 nrs=146.667e-3 sa=440e-9
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M185 n259 n335 VDD VDD pmos_6p0 m=1.0 w=3e-6 l=700e-9 nf=1.0 as=1.32e-12
+ ad=1.32e-12 ps=6.88e-6 pd=6.88e-6 nrd=146.667e-3 nrs=146.667e-3 sa=440e-9
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M186 n342 n335 VSS VSS nmos_6p0 m=1.0 w=3e-6 l=700e-9 nf=1.0 as=1.32e-12
+ ad=1.32e-12 ps=6.88e-6 pd=6.88e-6 nrd=146.667e-3 nrs=146.667e-3 sa=440e-9
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M187 n259 PD n342 VSS nmos_6p0 m=1.0 w=3e-6 l=700e-9 nf=1.0 as=1.32e-12
+ ad=1.32e-12 ps=6.88e-6 pd=6.88e-6 nrd=146.667e-3 nrs=146.667e-3 sa=440e-9
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M188 n348 n354 n335 VDD pmos_6p0 m=1.0 w=3e-6 l=700e-9 nf=1.0 as=1.32e-12
+ ad=1.32e-12 ps=6.88e-6 pd=6.88e-6 nrd=146.667e-3 nrs=146.667e-3 sa=440e-9
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M189 PU PD n335 VDD pmos_6p0 m=1.0 w=3e-6 l=700e-9 nf=1.0 as=1.32e-12
+ ad=1.32e-12 ps=6.88e-6 pd=6.88e-6 nrd=146.667e-3 nrs=146.667e-3 sa=440e-9
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M190 n354 PD VDD VDD pmos_6p0 m=1.0 w=3e-6 l=700e-9 nf=1.0 as=1.32e-12
+ ad=1.32e-12 ps=6.88e-6 pd=6.88e-6 nrd=146.667e-3 nrs=146.667e-3 sa=440e-9
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M191 n348 PU VDD VDD pmos_6p0 m=1.0 w=3e-6 l=700e-9 nf=1.0 as=1.32e-12
+ ad=1.32e-12 ps=6.88e-6 pd=6.88e-6 nrd=146.667e-3 nrs=146.667e-3 sa=440e-9
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M192 n348 PD n335 VSS nmos_6p0 m=1.0 w=1.5e-6 l=700e-9 nf=1.0 as=660e-15
+ ad=660e-15 ps=3.88e-6 pd=3.88e-6 nrd=293.333e-3 nrs=293.333e-3 sa=440e-9
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M193 PU n354 n335 VSS nmos_6p0 m=1.0 w=1.5e-6 l=700e-9 nf=1.0 as=660e-15
+ ad=660e-15 ps=3.88e-6 pd=3.88e-6 nrd=293.333e-3 nrs=293.333e-3 sa=440e-9
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M194 n354 PD VSS VSS nmos_6p0 m=1.0 w=1.5e-6 l=700e-9 nf=1.0 as=660e-15
+ ad=660e-15 ps=3.88e-6 pd=3.88e-6 nrd=293.333e-3 nrs=293.333e-3 sa=440e-9
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M195 n348 PU VSS VSS nmos_6p0 m=1.0 w=1.5e-6 l=700e-9 nf=1.0 as=660e-15
+ ad=660e-15 ps=3.88e-6 pd=3.88e-6 nrd=293.333e-3 nrs=293.333e-3 sa=440e-9
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
R196 n15 n357 $SUB=DVDD $[ppolyf_u] $W=800e-9 $L=23e-6 m=1.0 r=9.94533e3 par=1
R197 n357 n356 $SUB=DVDD $[ppolyf_u] $W=800e-9 $L=35.7e-6 m=1.0 r=15.3065e3 par=1
R198 n356 n355 $SUB=DVDD $[ppolyf_u] $W=800e-9 $L=35.7e-6 m=1.0 r=15.3065e3 par=1
R199 n355 n358 $SUB=DVDD $[ppolyf_u] $W=800e-9 $L=35.7e-6 m=1.0 r=15.3065e3 par=1
R200 n358 n363 $SUB=DVDD $[ppolyf_u] $W=800e-9 $L=35.7e-6 m=1.0 r=15.3065e3 par=1
R201 n363 n362 $SUB=DVDD $[ppolyf_u] $W=800e-9 $L=35.7e-6 m=1.0 r=15.3065e3 par=1
R202 n362 n359 $SUB=DVDD $[ppolyf_u] $W=800e-9 $L=35.7e-6 m=1.0 r=15.3065e3 par=1
R203 n359 n360 $SUB=DVDD $[ppolyf_u] $W=800e-9 $L=35.7e-6 m=1.0 r=15.3065e3 par=1
M204 n360 n276 DVSS DVSS nmos_6p0 m=1.0 w=1.5e-6 l=700e-9 nf=1.0 as=660e-15
+ ad=660e-15 ps=3.88e-6 pd=3.88e-6 nrd=293.333e-3 nrs=293.333e-3 sa=440e-9
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M205 n360 n260 DVDD DVDD pmos_6p0 m=1.0 w=3e-6 l=700e-9 nf=1.0 as=1.32e-12
+ ad=1.32e-12 ps=6.88e-6 pd=6.88e-6 nrd=146.667e-3 nrs=146.667e-3 sa=440e-9
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
D206 DVSS n15 np_6p0 m=2.0 AREA=20e-12 PJ=42e-6
D207 n15 DVDD pn_6p0 m=2.0 AREA=20e-12 PJ=42e-6
R208 PAD n15 $SUB=DVDD $[ppolyf_u] $W=2.5e-6 $L=2.8e-6 m=1.0 r=432.59 par=1
R209 PAD n15 $SUB=DVDD $[ppolyf_u] $W=2.5e-6 $L=2.8e-6 m=1.0 r=449.157 par=1
R210 PAD n15 $SUB=DVDD $[ppolyf_u] $W=2.5e-6 $L=2.8e-6 m=1.0 r=432.59 par=1
R211 PAD n15 $SUB=DVDD $[ppolyf_u] $W=2.5e-6 $L=2.8e-6 m=1.0 r=449.157 par=1
.ENDS
