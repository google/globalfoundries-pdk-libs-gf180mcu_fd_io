# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_io__fillnc
  CLASS PAD SPACER ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_fd_io__fillnc 0 0 ;
  SIZE 0.1 BY 350 ;
  SYMMETRY X Y R90 ;
  SITE GF_IO_Site ;
  PIN DVDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal3 ;
        RECT 0 334 0.1 341 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0 294 0.1 301 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0 278 0.1 285 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0 270 0.1 277 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0 262 0.1 269 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0 214 0.1 229 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0 206 0.1 213 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0 182 0.1 197 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0 166 0.1 181 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0 150 0.1 165 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0 134 0.1 149 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 0 334 0.1 341 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 0 294 0.1 301 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 0 278 0.1 285 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 0 270 0.1 277 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 0 262 0.1 269 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 0 214 0.1 229 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 0 206 0.1 213 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 0 182 0.1 197 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 0 166 0.1 181 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 0 150 0.1 165 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 0 134 0.1 149 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 0 334 0.1 341 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 0 294 0.1 301 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 0 278 0.1 285 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 0 270 0.1 277 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 0 262 0.1 269 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 0 214 0.1 229 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 0 206 0.1 213 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 0 182 0.1 197 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 0 166 0.1 181 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 0 150 0.1 165 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 0 134 0.1 149 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 0 118 0.1 125 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 0 118 0.1 125 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0 118 0.1 125 ;
    END
  END DVDD
  PIN DVSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal3 ;
        RECT 0 342 0.1 348.39 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0 326 0.1 333 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0 302 0.1 309 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0 286 0.1 293 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0 230 0.1 245 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0 198 0.1 205 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0 126 0.1 133 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0 102 0.1 117 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0 86 0.1 101 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 0 342 0.1 348.39 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 0 326 0.1 333 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 0 302 0.1 309 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 0 286 0.1 293 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 0 230 0.1 245 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 0 198 0.1 205 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 0 126 0.1 133 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 0 102 0.1 117 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 0 86 0.1 101 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 0 342 0.1 348.39 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 0 326 0.1 333 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 0 302 0.1 309 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 0 286 0.1 293 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 0 230 0.1 245 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 0 198 0.1 205 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 0 126 0.1 133 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 0 102 0.1 117 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 0 86 0.1 101 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 0 70 0.1 85 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 0 70 0.1 85 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0 70 0.1 85 ;
    END
  END DVSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal3 ;
        RECT 0 310 0.1 317 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 0 310 0.1 317 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 0 310 0.1 317 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 0 254 0.1 261 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 0 254 0.1 261 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0 254 0.1 261 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal3 ;
        RECT 0 318 0.1 325 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 0 318 0.1 325 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 0 318 0.1 325 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 0 246 0.1 253 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 0 246 0.1 253 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0 246 0.1 253 ;
    END
  END VSS
  OBS
    LAYER Metal1 ;
      RECT 0 0 0.1 350 ;
    LAYER Metal2 ;
      RECT 0 0 0.1 350 ;
    LAYER Metal3 ;
      RECT 0 341.28 0.1 341.72 ;
      RECT 0 165.28 0.1 165.72 ;
      RECT 0 245.28 0.1 245.72 ;
      RECT 0 125.28 0.1 125.72 ;
      RECT 0 253.28 0.1 253.72 ;
      RECT 0 277.28 0.1 277.72 ;
      RECT 0 309.28 0.1 309.72 ;
      RECT 0 133.28 0.1 133.72 ;
      RECT 0 269.28 0.1 269.72 ;
      RECT 0 229.28 0.1 229.72 ;
      RECT 0 348.67 0.1 350 ;
      RECT 0 293.28 0.1 293.72 ;
      RECT 0 317.28 0.1 317.72 ;
      RECT 0 285.28 0.1 285.72 ;
      RECT 0 213.28 0.1 213.72 ;
      RECT 0 261.28 0.1 261.72 ;
      RECT 0 101.28 0.1 101.72 ;
      RECT 0 205.28 0.1 205.72 ;
      RECT 0 333.28 0.1 333.72 ;
      RECT 0 197.28 0.1 197.72 ;
      RECT 0 181.28 0.1 181.72 ;
      RECT 0 301.28 0.1 301.72 ;
      RECT 0 149.28 0.1 149.72 ;
      RECT 0 0 0.1 69.72 ;
      RECT 0 85.28 0.1 85.72 ;
      RECT 0 117.28 0.1 117.72 ;
      RECT 0 325.28 0.1 325.72 ;
    LAYER Metal4 ;
      RECT 0 181.28 0.1 181.72 ;
      RECT 0 229.28 0.1 229.72 ;
      RECT 0 245.28 0.1 245.72 ;
      RECT 0 285.28 0.1 285.72 ;
      RECT 0 277.28 0.1 277.72 ;
      RECT 0 85.28 0.1 85.72 ;
      RECT 0 125.28 0.1 125.72 ;
      RECT 0 149.28 0.1 149.72 ;
      RECT 0 0 0.1 69.72 ;
      RECT 0 341.28 0.1 341.72 ;
      RECT 0 117.28 0.1 117.72 ;
      RECT 0 348.67 0.1 350 ;
      RECT 0 197.28 0.1 197.72 ;
      RECT 0 309.28 0.1 309.72 ;
      RECT 0 301.28 0.1 301.72 ;
      RECT 0 317.28 0.1 317.72 ;
      RECT 0 133.28 0.1 133.72 ;
      RECT 0 269.28 0.1 269.72 ;
      RECT 0 205.28 0.1 205.72 ;
      RECT 0 293.28 0.1 293.72 ;
      RECT 0 253.28 0.1 253.72 ;
      RECT 0 165.28 0.1 165.72 ;
      RECT 0 213.28 0.1 213.72 ;
      RECT 0 261.28 0.1 261.72 ;
      RECT 0 325.28 0.1 325.72 ;
      RECT 0 333.28 0.1 333.72 ;
      RECT 0 101.28 0.1 101.72 ;
    LAYER Metal5 ;
      RECT 0 125.28 0.1 125.72 ;
      RECT 0 165.28 0.1 165.72 ;
      RECT 0 333.28 0.1 333.72 ;
      RECT 0 285.28 0.1 285.72 ;
      RECT 0 309.28 0.1 309.72 ;
      RECT 0 133.28 0.1 133.72 ;
      RECT 0 85.28 0.1 85.72 ;
      RECT 0 149.28 0.1 149.72 ;
      RECT 0 348.67 0.1 350 ;
      RECT 0 229.28 0.1 229.72 ;
      RECT 0 197.28 0.1 197.72 ;
      RECT 0 317.28 0.1 317.72 ;
      RECT 0 269.28 0.1 269.72 ;
      RECT 0 181.28 0.1 181.72 ;
      RECT 0 101.28 0.1 101.72 ;
      RECT 0 261.28 0.1 261.72 ;
      RECT 0 0 0.1 69.72 ;
      RECT 0 245.28 0.1 245.72 ;
      RECT 0 253.28 0.1 253.72 ;
      RECT 0 205.28 0.1 205.72 ;
      RECT 0 213.28 0.1 213.72 ;
      RECT 0 277.28 0.1 277.72 ;
      RECT 0 117.28 0.1 117.72 ;
      RECT 0 293.28 0.1 293.72 ;
      RECT 0 325.28 0.1 325.72 ;
      RECT 0 341.28 0.1 341.72 ;
      RECT 0 301.28 0.1 301.72 ;
    LAYER Via1 ;
      RECT 0 0 0.1 350 ;
    LAYER Via2 ;
      RECT 0 0 0.1 350 ;
    LAYER Via3 ;
      RECT 0 0 0.1 350 ;
    LAYER Via4 ;
      RECT 0 0 0.1 350 ;
  END

END gf180mcu_fd_io__fillnc
